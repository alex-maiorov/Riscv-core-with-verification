// The actual core will be here